package <uvc_name>_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "<uvc_name>_config.svh"
  `include "<uvc_name>_seq_item.svh"
  `include "<uvc_name>_driver.svh"
  `include "<uvc_name>_monitor.svh"
  `include "<uvc_name>_seq_base.svh"
  `include "<uvc_name>_agent.svh"
endpackage:<uvc_name>_pkg
